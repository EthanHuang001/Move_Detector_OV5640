
`timescale 1ns / 1ns
module CMOS_OVxxxx_RGB640480
(
	//global clock 50MHz
	input			clk,			//50MHz
	input			rst_n,			//global reset
	
	//sdram1 control
	output			sdram1_clk,		//sdram clock
	output			sdram1_cke,		//sdram clock enable
	output			sdram1_cs_n,		//sdram chip select
	output			sdram1_we_n,		//sdram write enable
	output			sdram1_cas_n,	//sdram column address strobe
	output			sdram1_ras_n,	//sdram row address strobe
   //output	[1:0]	sdram1_dqm,		//sdram data enable
	output	[1:0]	sdram1_ba,		//sdram bank address
	output	[12:0]  sdram1_addr,		//sdram address
	inout	[15:0]	sdram1_data,		//sdram data
	
	//sdram2 control
	output			sdram2_clk,		//sdram clock
	output			sdram2_cke,		//sdram clock enable
	output			sdram2_cs_n,		//sdram chip select
	output			sdram2_we_n,		//sdram write enable
	output			sdram2_cas_n,	//sdram column address strobe
	output			sdram2_ras_n,	//sdram row address strobe
   //output	[1:0]	sdram2_dqm,		//sdram data enable
	output	[1:0]	sdram2_ba,		//sdram bank address
	output	[12:0]  sdram2_addr,		//sdram address
	inout	[15:0]	sdram2_data,		//sdram data
	
	//lcd port
//	output			lcd_dclk,		//lcd pixel clock			
	output			lcd_hs,			//lcd horizontal sync 
	output			lcd_vs,			//lcd vertical sync
//	output			lcd_sync,		//lcd sync
//	output			lcd_blank,		//lcd blank(L:blank)
//	output			lcd_de,			//lcd data enable
	output	[4:0]	lcd_red,		//lcd red data
	output	[5:0]	lcd_green,		//lcd green data
	output	[4:0]	lcd_blue,		//lcd blue data
   
   //gray_port
   output			gray_hs,			//gray horizontal sync 
	output			gray_vs,			//gray vertical sync
	output	[7:0]	gray_data,		//gray data

	//cmos interface
    //����ͷ�ӿ�
    input                 cam_pclk    ,  //cmos ��������ʱ��
	 output                cam_xclk    ,
    input                 cam_vsync   ,  //cmos ��ͬ���ź�
    input                 cam_href    ,  //cmos ��ͬ���ź�
    input        [7:0]    cam_data    ,  //cmos ����  
    output                cam_rst_n   ,  //cmos ��λ�źţ��͵�ƽ��Ч
    output                cam_pwdn    ,  //cmos ��Դ����ģʽѡ���ź�
    output                cam_scl     ,  //cmos SCCB_SCL��
    inout                 cam_sda       //cmos SCCB_SDA��
	

);


wire[15:0]                      vout_data;
assign lcd_red   = {vout_data[15:11]};
assign lcd_green = {vout_data[10:5]};
assign lcd_blue  = {vout_data[4:0]};

//---------------------------------------------
//system global clock control
wire	sys_rst_n;		//global reset
wire	clk_ref;		//sdram ctrl clock
wire	clk_refout;		//sdram clock output
wire	clk_vga;		//vga clock
//wire	clk_cmos;		//24MHz cmos clock
//wire	clk_48M;		//48MHz SignalTap II Clock


system_ctrl_pll	u_system_ctrl_pll
(
	.clk				(clk),			//global clock
	.rst_n				(rst_n),		//external reset
	
	.sys_rst_n			(sys_rst_n),	//global reset
	.clk_c0				(clk_ref),		//100MHz 
	.clk_c1				(clk_refout),	//100MHz -90deg
	.clk_c2				(clk_vga),		//25MHz
	.clk_c3				(cam_xclk)	//24MHz
);
//----------------------------------------------
//parameter define
parameter  SLAVE_ADDR = 7'h3c         ;  //OV5640��������ַ7'h3c
parameter  BIT_CTRL   = 1'b1          ;  //OV5640���ֽڵ�ַΪ16λ  0:8λ 1:16λ
parameter  CLK_FREQ   = 26'd25_000_000;  //i2c_driģ�������ʱ��Ƶ�� 25MHz
parameter  I2C_FREQ   = 18'd250_000   ;  //I2C��SCLʱ��Ƶ��,������400KHz
parameter  CMOS_H_PIXEL = 24'd640     ;  //CMOSˮƽ�������ظ���,��������SDRAM�����С
parameter  CMOS_V_PIXEL = 24'd480     ;  //CMOS��ֱ�������ظ���,��������SDRAM�����С
wire                  i2c_exec        ;  //I2C����ִ���ź�
wire   [23:0]         i2c_data        ;  //I2CҪ���õĵ�ַ������(��8λ��ַ,��8λ����)          
wire                  cam_init_done   ;  //����ͷ��ʼ�����
wire	    	      sdram_init_done;			//sdram init done
wire                  i2c_done        ;  //I2C�Ĵ�����������ź�
wire                  i2c_dri_clk     ;  //I2C����ʱ��
//��������ͷӲ����λ,�̶��ߵ�ƽ
assign  cam_rst_n = 1'b1;
//��Դ����ģʽѡ�� 0������ģʽ 1����Դ����ģʽ
assign  cam_pwdn = 1'b0;
 //I2C����ģ��
i2c_ov5640_rgb565_cfg 
   #(
     .CMOS_H_PIXEL  (CMOS_H_PIXEL),
     .CMOS_V_PIXEL  (CMOS_V_PIXEL)
    )
   u_i2c_cfg(
    .clk           (i2c_dri_clk),
    .rst_n         (rst_n),
    .i2c_done      (i2c_done),
    .i2c_exec      (i2c_exec),
    .i2c_data      (i2c_data),
    .init_done     (cam_init_done)
    );    

//I2C����ģ��
i2c_dri 
   #(
    .SLAVE_ADDR  (SLAVE_ADDR),               //��������
    .CLK_FREQ    (CLK_FREQ  ),              
    .I2C_FREQ    (I2C_FREQ  )                
    ) 
   u_i2c_dri(
    .clk         (clk_vga   ),//25M
    .rst_n       (rst_n     ),   
    //i2c interface
    .i2c_exec    (i2c_exec  ),   
    .bit_ctrl    (BIT_CTRL  ),   
    .i2c_rh_wl   (1'b0),                     //�̶�Ϊ0��ֻ�õ���IIC������д����   
    .i2c_addr    (i2c_data[23:8]),   
    .i2c_data_w  (i2c_data[7:0]),   
    .i2c_data_r  (),   
    .i2c_done    (i2c_done  ),   
    .scl         (cam_scl   ),   
    .sda         (cam_sda   ),   
    //user interface
    .dri_clk     (i2c_dri_clk)               //I2C����ʱ��
);
//CMOSͼ�����ݲɼ�ģ��
wire			cmos_frame_vsync;	//cmos frame data vsync valid signal
wire			cmos_frame_href;	//cmos frame data href vaild  signal
wire	[15:0]	cmos_frame_data;	//cmos frame data output: {cmos_data[7:0]<<8, cmos_data[7:0]}	
wire			cmos_frame_clken;	//cmos frame data output/capture enable clock
cmos_capture_data u_cmos_capture_data(
    .rst_n               (rst_n & cam_init_done), //ϵͳ��ʼ�����֮���ٿ�ʼ�ɼ����� 
    .cam_pclk            (cam_pclk),
    .cam_vsync           (!cam_vsync),
    .cam_href            (cam_href),
    .cam_data            (cam_data),         
    .cmos_frame_vsync    (cmos_frame_vsync),
    .cmos_frame_href     (cmos_frame_href),
    .cmos_frame_valid    (cmos_frame_clken),            //������Чʹ���ź�
    .cmos_frame_data     (cmos_frame_data)           //��Ч���� 
    );

//--------------------------------------------------------------------------------------
//--------------------------------------------------------------------------------------
//cmos video image capture

//wire	[7:0]	led_data = cmos_fps_rate;
wire        lcd_request             ;
//wire	[7:0]	led_data = LUT_INDEX;
//wire	[7:0]	led_data = i2c_rdata;

//********************************************
wire [15:0]  gray_sft; 
wire         sdr_rd; 
wire         gs_clken ;
wire         post_frame_vsync;
wire         post_frame_href;
wire [15:0]  post_img_data;
wire         post_frame_clken;
//-------------------------------------


//Sdram_Control_4Port module 	
//sdram write port1
wire			 sdr_wr1_clk	  = cam_pclk     ;	//Change with input signal											
wire	[7:0]  sdr_wr1_wrdata  = gray_sft[15:8];
wire			 sdr_wr1_wrreq   = gs_clken ;//gs_clken ;

//sdram read  port1
wire			 sdr_rd1_clk	  = cam_pclk ;	//Change with vga timing	
wire	[7:0]  sys_data_out1   ;
wire			 sys_rd1         = sdr_rd ;
wire         RD1_EMPTY;


//sdram write port2
wire			 sdr_wr2_clk	  =   cam_pclk;	//Change with input signal											
wire	[15:0] sdr_wr2_wrdata  =   post_img_data ;// {16{post_img_Bit}};//{data_diff,data_diff}; //sys_data_sim for test
wire			 sdr_wr2_wrreq   =   post_frame_clken;//sys_we_sim for test
//sdram read  port2
wire			 sdr_rd2_clk	=	clk_vga;	//Change with vga timing	
wire	[15:0] sys_data_out2;
wire			 sys_rd2       =  lcd_request;
wire         RD2_EMPTY;



Video_Image_Processor 
#(
	.IMG_HDISP(10'd640),	//640*48s0
	.IMG_VDISP(10'd480)
)
Video_Image_Processor_u0
(
	//global clock
	.clk				   	(cam_pclk),  			//cmos video pixel clock
	.rst_n					(sys_rst_n),			//global reset
	.cmos_frame_clken		(cmos_frame_clken), 	//Prepared Image data vsync valid signal
	.cmos_frame_vsync		(cmos_frame_vsync), 		//Prepared Image data href vaild  signal
	.cmos_frame_href		(cmos_frame_href ), 	//Prepared Image data output/capture enable clock
	.cmos_frame_data     (cmos_frame_data),			//Prepared Image brightness input
	//Image data has been processd
	.post_frame_vsync    (post_frame_vsync),
	.post_frame_href		(post_frame_href),		//Processed Image data href vaild  signal
	.post_frame_clken		(post_frame_clken),		//Processed Image data output/capture enable clock
	.post_img_data       (post_img_data),			//Processed Image brightness output
	.sys_data_out1       (sys_data_out1),
	.gs_clken            (gs_clken),
	.gray_sft            (gray_sft),
	.sdr_rd              (sdr_rd),
.gs_vsync(gs_vsync),
	//user interface
	.Sobel_Threshold     ( 8'd20 )		// 8'd10 ~8'd20
);
wire gs_vsync;
//wire sdram_init_done;
	/*Sdram_Control_4Port Sdram_Control_4Port(
		//	HOST Side
		.REF_CLK(clk_ref),
		.OUT_CLK(clk_refout),
		.RESET_N(sys_rst_n),	//��λ���룬�͵�ƽ��λ
		//.SDRAM_INIT_DONE(sdram_init_done),
		//	FIFO Write Side 1
		.WR1_DATA(sdr_wr1_wrdata),			//д��˿�1����������ˣ�16bit
		.WR1(sdr_wr1_wrreq),					//д��˿�1��дʹ�ܶˣ��ߵ�ƽд��
		.WR1_ADDR(0),			//д��˿�1��д��ʼ��ַ
		.WR1_MAX_ADDR(640*480-1),		//д��˿�1��д������ַ
		.WR1_LENGTH(256),			//һ����д�����ݳ���
		.WR1_LOAD(~sys_rst_n),			//д��˿�1�������󣬸ߵ�ƽ����д���ַ��fifo
		.WR1_CLK(sdr_wr1_clk),				//д��˿�1 fifoд��ʱ��
		.WR1_FULL(),			//д��˿�1 fifoд���ź�
		.WR1_USE(),				//д��˿�1 fifo�Ѿ�д������ݳ���

		//	FIFO Write Side 2
		.WR2_DATA(sdr_wr2_wrdata),			//д��˿�2����������ˣ�16bit
		.WR2(sdr_wr2_wrreq),					//д��˿�2��дʹ�ܶˣ��ߵ�ƽд��
		.WR2_ADDR(640*480),			//д��˿�2��д��ʼ��ַ
		.WR2_MAX_ADDR(640*480*2-1),		//д��˿�2��д������ַ
		.WR2_LENGTH(256),			//һ����д�����ݳ���
		.WR2_LOAD(~sys_rst_n),			//д��˿�2�������󣬸ߵ�ƽ����д���ַ��fifo
		.WR2_CLK(sdr_wr2_clk),				//д��˿�2 fifoд��ʱ��
		.WR2_FULL(),			//д��˿�2 fifoд���ź�
		.WR2_USE(),				//д��˿�2 fifo�Ѿ�д������ݳ���

		//	FIFO Read Side 1
		.RD1_DATA(sys_data_out1),			//�����˿�1����������ˣ�16bit
		.RD1(sys_rd1),					//�����˿�1�Ķ�ʹ�ܶˣ��ߵ�ƽ����
		.RD1_ADDR(0),			//�����˿�1�Ķ���ʼ��ַ
		.RD1_MAX_ADDR(640*480-1),		//�����˿�1�Ķ�������ַ
		.RD1_LENGTH(128),			//һ���Զ������ݳ���
		.RD1_LOAD(~sys_rst_n),			//�����˿�1 �������󣬸ߵ�ƽ���������ַ��fifo
		.RD1_CLK(sdr_rd1_clk),				//�����˿�1 fifo��ȡʱ��
		.RD1_EMPTY(RD1_EMPTY),			//�����˿�1 fifo�����ź�
		.RD1_USE(),				//�����˿�1 fifo�Ѿ������Զ�ȡ�����ݳ���

		//	FIFO Read Side 2
		.RD2_DATA(sys_data_out2),			//�����˿�2����������ˣ�16bit
		.RD2(sys_rd2),					//�����˿�2�Ķ�ʹ�ܶˣ��ߵ�ƽ����
		.RD2_ADDR(640*480),			//�����˿�2�Ķ���ʼ��ַ
		.RD2_MAX_ADDR(640*480*2-1),		//�����˿�2�Ķ�������ַ
		.RD2_LENGTH(128),			//һ���Զ������ݳ���
		.RD2_LOAD(~sys_rst_n),			//�����˿�2�������󣬸ߵ�ƽ���������ַ��fifo
		.RD2_CLK(sdr_rd2_clk),				//�����˿�2 fifo��ȡʱ��
		.RD2_EMPTY(RD2_EMPTY),			//�����˿�2 fifo�����ź�
		.RD2_USE(),				//�����˿�2 fifo�Ѿ������Զ�ȡ�����ݳ���

		//	SDRAM Side
		
		.SA(sdram_addr),		//SDRAM ��ַ�ߣ�
		.BA(sdram_ba),		//SDRAM bank��ַ��
		.CS_N(sdram_cs_n),		//SDRAM Ƭѡ�ź�
		.CKE(sdram_cke),		//SDRAM ʱ��ʹ��
		.RAS_N(sdram_ras_n),	//SDRAM ��ѡ���ź�
		.CAS_N(sdram_cas_n),	//SDRAM ��ѡ���ź�
		.WE_N(sdram_we_n),		//SDRAM д�����ź�
		.DQ(sdram_data),		//SDRAM ˫����������
		.SDR_CLK(sdram_clk),
		.DQM(sdram_dqm),		//SDRAM �������߸ߵ��ֽ������ź�
		.Sdram_Init_Done(sdram_init_done)
	);
*/
wire sdram1_init_done;
wire sdram2_init_done;
sdram_top   sdram1_top_inst(

    .sys_clk            (clk_ref    ),  //sdram �������ο�ʱ��
    .clk_out            (clk_refout ),  //�����������λƫ��ʱ��
    .sys_rst_n          (sys_rst_n         ),  //ϵͳ��λ
//�û�д�˿�
    .wr_fifo_wr_clk     (sdr_wr1_clk    ),  //д�˿�FIFO: дʱ��
    .wr_fifo_wr_req     (sdr_wr1_wrreq  ),  //д�˿�FIFO: дʹ��
    .wr_fifo_wr_data    (sdr_wr1_wrdata ),  //д�˿�FIFO: д����
    .sdram_wr_b_addr    (24'd0          ),  //дSDRAM����ʼ��ַ
    .sdram_wr_e_addr    (640*480        ),  //дSDRAM�Ľ�����ַ
    .wr_burst_len       (10'd512        ),  //дSDRAMʱ������ͻ�����ȁ8�2�8�2
    .wr_rst             (~rst_n         ),  //д�˿ڸ�λ: ��λд��ַ,���дFIFO
//�û����˿�
    .rd_fifo_rd_clk     (sdr_rd1_clk    ),  //���˿�FIFO: ��ʱ��
    .rd_fifo_rd_req     (sys_rd1        ),  //���˿�FIFO: ��ʹ��
    .rd_fifo_rd_data    (sys_data_out1  ),  //���˿�FIFO: ������
    .sdram_rd_b_addr    (24'd0          ),  //��SDRAM����ʼ��ַ
    .sdram_rd_e_addr    (640*480        ),  //��SDRAM�Ľ�����ַ
    .rd_burst_len       (10'd512        ),  //��SDRAM�ж�����ʱ��ͻ������
    .rd_rst             (~sys_rst_n     ),  //���˿ڸ�λ: ��λ����ַ,��ն�FIFO
	.rdempty            (RD1_EMPTY      ),   //�����ź�
//�û����ƶ˿�
    .read_valid         (1'b1           ),  //SDRAM ��ʹ��
    .pingpang_en        (1'b1           ),  //SDRAM ƹ�Ҳ���ʹ��
    .init_end           (sdram1_init_done),  //SDRAM ��ʼ����ɱ�־
//SDRAM оƬ�ӿ�
    .sdram_clk          (sdram1_clk      ),  //SDRAM оƬʱ��
    .sdram_cke          (sdram1_cke      ),  //SDRAM ʱ����Ч
    .sdram_cs_n         (sdram1_cs_n     ),  //SDRAM Ƭѡ
    .sdram_ras_n        (sdram1_ras_n    ),  //SDRAM ����Ч
    .sdram_cas_n        (sdram1_cas_n    ),  //SDRAM ����Ч
    .sdram_we_n         (sdram1_we_n     ),  //SDRAM д��Ч
    .sdram_ba           (sdram1_ba       ),  //SDRAM Bank��ַ
    .sdram_addr         (sdram1_addr     ),  //SDRAM ��/�е�ַ
    .sdram_dq           (sdram1_data      )  //SDRAM ����


);


sdram_top   sdram2_top_inst(

    .sys_clk            (clk_ref    ),  //sdram �������ο�ʱ��
    .clk_out            (clk_refout ),  //�����������λƫ��ʱ��
    .sys_rst_n          (sys_rst_n         ),  //ϵͳ��λ
//�û�д�˿�
    .wr_fifo_wr_clk     (sdr_wr2_clk    ),  //д�˿�FIFO: дʱ��
    .wr_fifo_wr_req     (sdr_wr2_wrreq  ),  //д�˿�FIFO: дʹ��
    .wr_fifo_wr_data    (sdr_wr2_wrdata ),  //д�˿�FIFO: д����
    .sdram_wr_b_addr    (24'd0          ),  //дSDRAM����ʼ��ַ
    .sdram_wr_e_addr    (640*480        ),  //дSDRAM�Ľ�����ַ
    .wr_burst_len       (10'd512        ),  //дSDRAMʱ������ͻ�����ȁ8�2�8�2
    .wr_rst             (~sys_rst_n     ),  //д�˿ڸ�λ: ��λд��ַ,���дFIFO
//�û����˿�
    .rd_fifo_rd_clk     (sdr_rd2_clk    ),  //���˿�FIFO: ��ʱ��
    .rd_fifo_rd_req     (sys_rd2        ),  //���˿�FIFO: ��ʹ��
    .rd_fifo_rd_data    (sys_data_out2  ),  //���˿�FIFO: ������
    .sdram_rd_b_addr    (24'd0          ),  //��SDRAM����ʼ��ַ
    .sdram_rd_e_addr    (640*480        ),  //��SDRAM�Ľ�����ַ
    .rd_burst_len       (10'd512        ),  //��SDRAM�ж�����ʱ��ͻ������
    .rd_rst             (~sys_rst_n     ),  //���˿ڸ�λ: ��λ����ַ,��ն�FIFO
	.rdempty            (RD2_EMPTY      ),   //�����ź�
//�û����ƶ˿�
    .read_valid         (1'b1           ),  //SDRAM ��ʹ��
    .pingpang_en        (1'b1           ),  //SDRAM ƹ�Ҳ���ʹ��
    .init_end           (sdram2_init_done),  //SDRAM ��ʼ����ɱ�־
//SDRAM оƬ�ӿ�
    .sdram_clk          (sdram2_clk      ),  //SDRAM оƬʱ��
    .sdram_cke          (sdram2_cke      ),  //SDRAM ʱ����Ч
    .sdram_cs_n         (sdram2_cs_n     ),  //SDRAM Ƭѡ
    .sdram_ras_n        (sdram2_ras_n    ),  //SDRAM ����Ч
    .sdram_cas_n        (sdram2_cas_n    ),  //SDRAM ����Ч
    .sdram_we_n         (sdram2_we_n     ),  //SDRAM д��Ч
    .sdram_ba           (sdram2_ba       ),  //SDRAM Bank��ַ
    .sdram_addr         (sdram2_addr     ),  //SDRAM ��/�е�ַ
    .sdram_dq           (sdram2_data      )  //SDRAM ����


);
//-------------------------------------
//LCD driver timing
lcd_driver u_lcd_driver
(
	//global clock
	.clk			(clk_vga),		
	.rst_n			(sys_rst_n), 
	 
	 //lcd interface
	.lcd_dclk		(),
	.lcd_blank		(),//lcd_blank
	.lcd_sync		(),		    	
	.lcd_hs			(lcd_hs),		
	.lcd_vs			(lcd_vs),
	.lcd_en			(),		
	.lcd_rgb		(vout_data),

	
	//user interface
	.lcd_request	(lcd_request),
	.lcd_data		(sys_data_out2),	
	.lcd_xpos		(),	
	.lcd_ypos		()
);
//GRAY driver timing
lcd_driver u_gray_driver
(
	//global clock
	.clk			(clk_vga),		
	.rst_n			(sys_rst_n), 
	 
	 //lcd interface
	.lcd_dclk		(),
	.lcd_blank		(),//lcd_blank
	.lcd_sync		(),		    	
	.lcd_hs			(gray_hs),		
	.lcd_vs			(gray_vs),
	.lcd_en			(),		
	.lcd_rgb		(gray_data),

	
	//user interface
	.lcd_request	(),
	.lcd_data		(sys_data_out1),	
	.lcd_xpos		(),	
	.lcd_ypos		()
);

endmodule
